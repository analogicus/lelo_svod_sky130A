*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_EXSC_lpe.spi
#else
.include ../../../work/xsch/LELO_EXSC.spice
#endif
.include ../../../design/1812PS.lib
.include ../../../design/XGL6030.lib
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  0 dc 40m
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.OPTIONS SAVECURRENTS
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.nodeset v(xdut.vddcs) = 0.6
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


tran 100n 1000u



write
quit


.endc

.end
