*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_EXSC_lpe.spi
#else
.include ../../../work/xsch/LELO_EXSC.spice
#endif
.include ../../../design/1812PS.lib
.include ../../../design/2014VS.lib
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  VSS dc 10m
VSS  VSS  0   dc 0
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.OPTIONS SAVECURRENTS
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


tran 500n 500u
let VDS3 = V(VDD)-V(xdut.VP1)
let VDS4 = V(xdut.VP1)-V(xdut.VP2)
let VDS5 = V(xdut.VP2)-V(xdut.VP3)
let VDS6 = V(xdut.VP3)-V(xdut.VP4)
let VDS7 = V(xdut.VP4)-V(xdut.vddcs)
save VDS3
save VDS4
save VDS5
save VDS6
save VDS7

write
quit


.endc

.end
