*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_CAP_lpe.spi
#else
.include ../../../work/xsch/LELO_CAP.spice
#endif
.include "/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt.pm3.spice"

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param freq = 1Meg
.csparam freq = {freq}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
IAC  VDD  VSS  dc 0 ac 1

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black

ac lin 10 1Meg 10Meg
* ac current source
echo impedance V/I:
*current in IAC normalized to 1 yields v(N4,N3)/1
print v(VDD,VSS)
echo conductance I/V = 1/R  + jwC
print 1/v(VDD,VSS)
echo capacitance
print imag(1/v(VDD,VSS))/2/PI/freq


.endc

.end
