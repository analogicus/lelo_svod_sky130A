*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_ONESHOT_VC_lpe.spi
#else
.include ../../../work/xsch/LELO_ONESHOT_VC.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p



*-----------------------------------------------------------------
* FORCE
*(0 0 10u 0.18 20u 0.36 30u 0.54 40u 0.72 50u 0.9 60u 1.08 70u 1.26 80u 1.44 90u 1.62 100u 1.8)
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS  dc 1.8
VC   VC   VSS  pwl 0 0 10u 0.18 20u 0.36 30u 0.54 40u 0.72 50u 0.9 60u 1.08 70u 1.26 80u 1.44 90u 1.62 100u 1.8
VIN   IN   VSS  PULSE(1.8 0 1n 1n 1n 5u 10u)
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 100n 110u
write
quit


.endc

.end
