*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_EXSC_lpe.spi
#else
.include ../../../work/xsch/LELO_EXSC.spice
#endif
.include ../../../work/xsch/1812PS.lib
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  VSS dc 4.5m
VSS  VSS  0   dc 0
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


tran 500n 1500u
let VG1_1 = V(xdut.VG1)
let VG2_1 = V(xdut.VG1)
save VG1
save VG2

write
quit


.endc

.end
