*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_BOOST_STEADY_STATE_lpe.spi
#else
.include ../../../work/xsch/LELO_BOOST_STEADY_STATE.spice
#endif
.include ../../../design/1812PS.lib
.include ../../../design/XGL6030.lib
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-5

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  0 dc 40m
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.OPTIONS SAVECURRENTS
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.nodeset v(xdut.teg) = 0.02
.nodeset v(xdut.vddc) = 1.8
.nodeset v(xdut.vc) = 0.65
.nodeset v(xdut.vc2) = 0.9

.control
set num_threads=8
set color0=white
set color1=black
unset askquit


tran 100n 100u



write
quit


.endc

.end
