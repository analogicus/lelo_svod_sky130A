*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_EXSC_lpe.spi
#else
.include ../../../work/xsch/LELO_EXSC.spice
#endif
.include ../../../design/1812PS.lib
.include ../../../design/XGL6030.lib
*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  0 dc 30m
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save @l.xdut.x7.x1.l1[i]
.save v(xdut.TEG)
.save v(xdut.VDDCS)
.save v(xdut.V1)
.save v(xdut.VHSS1)
.save v(xdut.VLSS)
.save v(xdut.vc)
.save v(xdut.x3.vg1)
.save v(xdut.x3.net3)
.save v(xdut.vdd_neg)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------

.nodeset v(xdut.teg) = 0.02
.nodeset v(xdut.VDDCS) = 0

.control
set num_threads=8
set color0=white
set color1=black
unset askquit


tran 100n 20000u



write
quit


.endc

.end
